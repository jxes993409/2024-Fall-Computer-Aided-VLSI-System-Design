// list all paths to your design files
`include "../01_RTL/core.v"
`include "../01_RTL/odd_even_sort.v"
`include "../01_RTL/divider.v"